module and12(input a,b, output out);

assign out = a&b;

endmodule
