`timescale 1ns/1ps
module CounterC (input clk,P,F,output [3:0] out_count);

reg[3:0]counter = 0;

always@(posedge clk)
begin
if (P == 1) begin
 if ( counter % 2 == 0) counter<=counter + 1; //set odd
 else if (F == 1) counter <= counter + 2;
 else counter <= counter - 2;
 end
else begin
if ( counter % 2 == 1) counter<=counter + 1; //set even
 else if (F == 1) counter <= counter + 2;
 else counter <= counter - 2;
end

end

endmodule
